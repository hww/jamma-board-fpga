library verilog;
use verilog.vl_types.all;
entity frontsextractor_6 is
    port(
        \P_c[13]\       : in     vl_logic;
        nreset_c_2      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i       : in     vl_logic;
        risea           : out    vl_logic
    );
end frontsextractor_6;
