library verilog;
use verilog.vl_types.all;
entity myfrontextractor_2 is
    port(
        \P_c[3]\        : in     vl_logic;
        nreset_c_0      : in     vl_logic;
        nreset_c_1      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i_0     : in     vl_logic;
        risea_n         : out    vl_logic
    );
end myfrontextractor_2;
