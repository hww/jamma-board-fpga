library verilog;
use verilog.vl_types.all;
entity frontsextractor is
    port(
        n_1097          : in     vl_logic;
        nreset_c_0      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i_0     : in     vl_logic;
        risea           : out    vl_logic
    );
end frontsextractor;
