library verilog;
use verilog.vl_types.all;
entity crt_measure_test is
end crt_measure_test;
