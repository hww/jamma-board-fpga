library verilog;
use verilog.vl_types.all;
entity mydffe2 is
    port(
        da_c            : in     vl_logic_vector(1 downto 0);
        dd_in_4         : in     vl_logic;
        dd_in_3         : in     vl_logic;
        dd_in_1         : in     vl_logic;
        dd_in_6         : in     vl_logic;
        dd_in_5         : in     vl_logic;
        dd_in_0         : in     vl_logic;
        key0            : out    vl_logic;
        nreset_c_3      : in     vl_logic;
        ndiow_c         : in     vl_logic;
        bdevice         : in     vl_logic;
        y_11            : in     vl_logic;
        cmd6n_0         : in     vl_logic;
        y_29            : in     vl_logic
    );
end mydffe2;
