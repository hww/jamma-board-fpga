library verilog;
use verilog.vl_types.all;
entity frontsextractor_4 is
    port(
        \P_c[11]\       : in     vl_logic;
        ndior_c_i       : in     vl_logic;
        nreset_c_1      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i_0     : in     vl_logic;
        risea           : out    vl_logic
    );
end frontsextractor_4;
