library verilog;
use verilog.vl_types.all;
entity frontsextractor_2 is
    port(
        nreset_c_0      : in     vl_logic;
        n_1069          : in     vl_logic;
        nreset_c_1      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i_0     : in     vl_logic;
        risea           : out    vl_logic
    );
end frontsextractor_2;
