library verilog;
use verilog.vl_types.all;
entity crt_top is
end crt_top;
