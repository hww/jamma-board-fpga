library verilog;
use verilog.vl_types.all;
entity frontsextractor_1 is
    port(
        n_1083          : in     vl_logic;
        nreset_c_0      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i_0     : in     vl_logic;
        riseb_n         : out    vl_logic
    );
end frontsextractor_1;
