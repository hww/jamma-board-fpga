library verilog;
use verilog.vl_types.all;
entity jamma is
    port(
        coincounter_c   : out    vl_logic_vector(2 downto 1);
        coinlockout_c   : out    vl_logic_vector(2 downto 1);
        dd_in           : in     vl_logic_vector(7 downto 0);
        bcounter        : out    vl_logic_vector(3 downto 0);
        da_c            : in     vl_logic_vector(2 downto 0);
        noice_1         : out    vl_logic;
        noice_2         : out    vl_logic;
        noice_15        : out    vl_logic;
        p_c_22          : in     vl_logic;
        p_c_12          : in     vl_logic;
        p_c_17          : in     vl_logic;
        p_c_7           : in     vl_logic;
        p_c_27          : in     vl_logic;
        p_c_24          : in     vl_logic;
        p_c_14          : in     vl_logic;
        p_c_28          : in     vl_logic;
        p_c_26          : in     vl_logic;
        p_c_25          : in     vl_logic;
        p_c_18          : in     vl_logic;
        p_c_8           : in     vl_logic;
        p_c_3           : in     vl_logic;
        p_c_16          : in     vl_logic;
        p_c_6           : in     vl_logic;
        p_c_1           : in     vl_logic;
        p_c_23          : in     vl_logic;
        p_c_13          : in     vl_logic;
        p_c_21          : in     vl_logic;
        p_c_11          : in     vl_logic;
        p_c_20          : in     vl_logic;
        p_c_10          : in     vl_logic;
        p_c_5           : in     vl_logic;
        p_c_0           : in     vl_logic;
        datainput_2     : out    vl_logic;
        datainput_0     : out    vl_logic;
        datainput_5     : out    vl_logic;
        datainput_4     : out    vl_logic;
        n_163           : in     vl_logic;
        ndior_c_i_0_0   : in     vl_logic;
        ndior_c_i       : in     vl_logic;
        clk_c           : in     vl_logic;
        ndiow_c         : in     vl_logic;
        y_3             : in     vl_logic;
        read            : out    vl_logic;
        ndior_c_i_0     : in     vl_logic;
        n_98            : out    vl_logic;
        n_105           : out    vl_logic;
        n_276           : in     vl_logic;
        n_110           : out    vl_logic;
        o1              : out    vl_logic;
        y_22            : out    vl_logic;
        y_27            : out    vl_logic;
        y_30            : out    vl_logic;
        y_33            : out    vl_logic;
        y_34            : out    vl_logic;
        nreset_c        : in     vl_logic;
        ndior_c         : in     vl_logic;
        ncs1_c          : in     vl_logic;
        ncs0_c          : in     vl_logic;
        acces           : out    vl_logic
    );
end jamma;
