library verilog;
use verilog.vl_types.all;
entity frontsextractor_3 is
    port(
        n_903           : in     vl_logic;
        nreset_c_1      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i_0     : in     vl_logic;
        riseb_n         : out    vl_logic
    );
end frontsextractor_3;
