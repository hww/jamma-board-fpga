library verilog;
use verilog.vl_types.all;
entity frontsextractor_7 is
    port(
        \P_c[14]\       : in     vl_logic;
        nreset_c_2      : in     vl_logic;
        clk_c           : in     vl_logic;
        ndior_c_i       : in     vl_logic;
        riseb_n         : out    vl_logic
    );
end frontsextractor_7;
